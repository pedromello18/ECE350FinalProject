module reg64(data_out, data_in, clk, writeEnable, reset);
    input [63:0] data_in;
    input clk, writeEnable, reset;

    output [63:0] data_out;

    dffe_ref BIT0(data_out[0], data_in[0], clk, writeEnable, reset);
    dffe_ref BIT1(data_out[1], data_in[1], clk, writeEnable, reset);
    dffe_ref BIT2(data_out[2], data_in[2], clk, writeEnable, reset);
    dffe_ref BIT3(data_out[3], data_in[3], clk, writeEnable, reset);
    dffe_ref BIT4(data_out[4], data_in[4], clk, writeEnable, reset);
    dffe_ref BIT5(data_out[5], data_in[5], clk, writeEnable, reset);
    dffe_ref BIT6(data_out[6], data_in[6], clk, writeEnable, reset);
    dffe_ref BIT7(data_out[7], data_in[7], clk, writeEnable, reset);
    dffe_ref BIT8(data_out[8], data_in[8], clk, writeEnable, reset);
    dffe_ref BIT9(data_out[9], data_in[9], clk, writeEnable, reset);
    dffe_ref BIT10(data_out[10], data_in[10], clk, writeEnable, reset);
    dffe_ref BIT11(data_out[11], data_in[11], clk, writeEnable, reset);
    dffe_ref BIT12(data_out[12], data_in[12], clk, writeEnable, reset);
    dffe_ref BIT13(data_out[13], data_in[13], clk, writeEnable, reset);
    dffe_ref BIT14(data_out[14], data_in[14], clk, writeEnable, reset);
    dffe_ref BIT15(data_out[15], data_in[15], clk, writeEnable, reset);
    dffe_ref BIT16(data_out[16], data_in[16], clk, writeEnable, reset);
    dffe_ref BIT17(data_out[17], data_in[17], clk, writeEnable, reset);
    dffe_ref BIT18(data_out[18], data_in[18], clk, writeEnable, reset);
    dffe_ref BIT19(data_out[19], data_in[19], clk, writeEnable, reset);
    dffe_ref BIT20(data_out[20], data_in[20], clk, writeEnable, reset);
    dffe_ref BIT21(data_out[21], data_in[21], clk, writeEnable, reset);
    dffe_ref BIT22(data_out[22], data_in[22], clk, writeEnable, reset);
    dffe_ref BIT23(data_out[23], data_in[23], clk, writeEnable, reset);
    dffe_ref BIT24(data_out[24], data_in[24], clk, writeEnable, reset);
    dffe_ref BIT25(data_out[25], data_in[25], clk, writeEnable, reset);
    dffe_ref BIT26(data_out[26], data_in[26], clk, writeEnable, reset);
    dffe_ref BIT27(data_out[27], data_in[27], clk, writeEnable, reset);
    dffe_ref BIT28(data_out[28], data_in[28], clk, writeEnable, reset);
    dffe_ref BIT29(data_out[29], data_in[29], clk, writeEnable, reset);
    dffe_ref BIT30(data_out[30], data_in[30], clk, writeEnable, reset);
    dffe_ref BIT31(data_out[31], data_in[31], clk, writeEnable, reset);
    dffe_ref BIT32(data_out[32], data_in[32], clk, writeEnable, reset);
    dffe_ref BIT33(data_out[33], data_in[33], clk, writeEnable, reset);
    dffe_ref BIT34(data_out[34], data_in[34], clk, writeEnable, reset);
    dffe_ref BIT35(data_out[35], data_in[35], clk, writeEnable, reset);
    dffe_ref BIT36(data_out[36], data_in[36], clk, writeEnable, reset);
    dffe_ref BIT37(data_out[37], data_in[37], clk, writeEnable, reset);
    dffe_ref BIT38(data_out[38], data_in[38], clk, writeEnable, reset);
    dffe_ref BIT39(data_out[39], data_in[39], clk, writeEnable, reset);
    dffe_ref BIT40(data_out[40], data_in[40], clk, writeEnable, reset);
    dffe_ref BIT41(data_out[41], data_in[41], clk, writeEnable, reset);
    dffe_ref BIT42(data_out[42], data_in[42], clk, writeEnable, reset);
    dffe_ref BIT43(data_out[43], data_in[43], clk, writeEnable, reset);
    dffe_ref BIT44(data_out[44], data_in[44], clk, writeEnable, reset);
    dffe_ref BIT45(data_out[45], data_in[45], clk, writeEnable, reset);
    dffe_ref BIT46(data_out[46], data_in[46], clk, writeEnable, reset);
    dffe_ref BIT47(data_out[47], data_in[47], clk, writeEnable, reset);
    dffe_ref BIT48(data_out[48], data_in[48], clk, writeEnable, reset);
    dffe_ref BIT49(data_out[49], data_in[49], clk, writeEnable, reset);
    dffe_ref BIT50(data_out[50], data_in[50], clk, writeEnable, reset);
    dffe_ref BIT51(data_out[51], data_in[51], clk, writeEnable, reset);
    dffe_ref BIT52(data_out[52], data_in[52], clk, writeEnable, reset);
    dffe_ref BIT53(data_out[53], data_in[53], clk, writeEnable, reset);
    dffe_ref BIT54(data_out[54], data_in[54], clk, writeEnable, reset);
    dffe_ref BIT55(data_out[55], data_in[55], clk, writeEnable, reset);
    dffe_ref BIT56(data_out[56], data_in[56], clk, writeEnable, reset);
    dffe_ref BIT57(data_out[57], data_in[57], clk, writeEnable, reset);
    dffe_ref BIT58(data_out[58], data_in[58], clk, writeEnable, reset);
    dffe_ref BIT59(data_out[59], data_in[59], clk, writeEnable, reset);
    dffe_ref BIT60(data_out[60], data_in[60], clk, writeEnable, reset);
    dffe_ref BIT61(data_out[61], data_in[61], clk, writeEnable, reset);
    dffe_ref BIT62(data_out[62], data_in[62], clk, writeEnable, reset);
    dffe_ref BIT63(data_out[63], data_in[63], clk, writeEnable, reset);

endmodule