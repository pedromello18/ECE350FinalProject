module ars_2(out, s, A);
    input s;
    input [64:0] A;
    output [64:0] out;

    mux_2 BIT0(out[0], s, A[0], A[2]);
    mux_2 BIT1(out[1], s, A[1], A[3]);
    mux_2 BIT2(out[2], s, A[2], A[4]);
    mux_2 BIT3(out[3], s, A[3], A[5]);
    mux_2 BIT4(out[4], s, A[4], A[6]);
    mux_2 BIT5(out[5], s, A[5], A[7]);
    mux_2 BIT6(out[6], s, A[6], A[8]);
    mux_2 BIT7(out[7], s, A[7], A[9]);
    mux_2 BIT8(out[8], s, A[8], A[10]);
    mux_2 BIT9(out[9], s, A[9], A[11]);
    mux_2 BIT10(out[10], s, A[10], A[12]);
    mux_2 BIT11(out[11], s, A[11], A[13]);
    mux_2 BIT12(out[12], s, A[12], A[14]);
    mux_2 BIT13(out[13], s, A[13], A[15]);
    mux_2 BIT14(out[14], s, A[14], A[16]);
    mux_2 BIT15(out[15], s, A[15], A[17]);
    mux_2 BIT16(out[16], s, A[16], A[18]);
    mux_2 BIT17(out[17], s, A[17], A[19]);
    mux_2 BIT18(out[18], s, A[18], A[20]);
    mux_2 BIT19(out[19], s, A[19], A[21]);
    mux_2 BIT20(out[20], s, A[20], A[22]);
    mux_2 BIT21(out[21], s, A[21], A[23]);
    mux_2 BIT22(out[22], s, A[22], A[24]);
    mux_2 BIT23(out[23], s, A[23], A[25]);
    mux_2 BIT24(out[24], s, A[24], A[26]);
    mux_2 BIT25(out[25], s, A[25], A[27]);
    mux_2 BIT26(out[26], s, A[26], A[28]);
    mux_2 BIT27(out[27], s, A[27], A[29]);
    mux_2 BIT28(out[28], s, A[28], A[30]);
    mux_2 BIT29(out[29], s, A[29], A[31]);
    mux_2 BIT30(out[30], s, A[30], A[32]);
    mux_2 BIT31(out[31], s, A[31], A[33]);
    mux_2 BIT32(out[32], s, A[32], A[34]);
    mux_2 BIT33(out[33], s, A[33], A[35]);
    mux_2 BIT34(out[34], s, A[34], A[36]);
    mux_2 BIT35(out[35], s, A[35], A[37]);
    mux_2 BIT36(out[36], s, A[36], A[38]);
    mux_2 BIT37(out[37], s, A[37], A[39]);
    mux_2 BIT38(out[38], s, A[38], A[40]);
    mux_2 BIT39(out[39], s, A[39], A[41]);
    mux_2 BIT40(out[40], s, A[40], A[42]);
    mux_2 BIT41(out[41], s, A[41], A[43]);
    mux_2 BIT42(out[42], s, A[42], A[44]);
    mux_2 BIT43(out[43], s, A[43], A[45]);
    mux_2 BIT44(out[44], s, A[44], A[46]);
    mux_2 BIT45(out[45], s, A[45], A[47]);
    mux_2 BIT46(out[46], s, A[46], A[48]);
    mux_2 BIT47(out[47], s, A[47], A[49]);
    mux_2 BIT48(out[48], s, A[48], A[50]);
    mux_2 BIT49(out[49], s, A[49], A[51]);
    mux_2 BIT50(out[50], s, A[50], A[52]);
    mux_2 BIT51(out[51], s, A[51], A[53]);
    mux_2 BIT52(out[52], s, A[52], A[54]);
    mux_2 BIT53(out[53], s, A[53], A[55]);
    mux_2 BIT54(out[54], s, A[54], A[56]);
    mux_2 BIT55(out[55], s, A[55], A[57]);
    mux_2 BIT56(out[56], s, A[56], A[58]);
    mux_2 BIT57(out[57], s, A[57], A[59]);
    mux_2 BIT58(out[58], s, A[58], A[60]);
    mux_2 BIT59(out[59], s, A[59], A[61]);
    mux_2 BIT60(out[60], s, A[60], A[62]);
    mux_2 BIT61(out[61], s, A[61], A[63]);
    mux_2 BIT62(out[62], s, A[62], A[64]);
    mux_2 BIT63(out[63], s, A[63], A[64]);
    mux_2 BIT64(out[64], s, A[64], A[64]);

endmodule